`timescale 1ns / 1ps//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 	 Alejandro Mora\Stiven Sanchez\Jorge Sequeira
// 
// Create Date:    01:53:12 01/05/2014 
// Design Name: 
// Module Name:    DECO_REF_POT
// Project Name: 	 Control Servo	
// Target Devices: 
// Tool versions: 
// Description: Decodificador que ecala el valor de REF a los valores correspondientes de POT
//////////////////////////////////////////////////////////////////////////////////
module DECO_REF_POT(IN,OUT);
	input [8:0] IN;
	output reg [7:0] OUT;
	
	always@(IN)
		case(IN)
			9'd20:OUT=8'b01110001;
			9'd21:OUT=8'b01110001;
			9'd22:OUT=8'b01110000;
			9'd23:OUT=8'b01101111;
			9'd24:OUT=8'b01101110;
			9'd25:OUT=8'b01101110;
			9'd26:OUT=8'b01101101;
			9'd27:OUT=8'b01101100;
			9'd28:OUT=8'b01101100;
			9'd29:OUT=8'b01101011;
			9'd30:OUT=8'b01101010;
			9'd31:OUT=8'b01101001;	
			9'd32:OUT=8'b01101001;
			9'd33:OUT=8'b01101000;
			9'd34:OUT=8'b01100111;
			9'd35:OUT=8'b01100111;
			9'd36:OUT=8'b01100110;
			9'd37:OUT=8'b01100101;
			9'd38:OUT=8'b01100100;
			9'd39:OUT=8'b01100100;
			9'd40:OUT=8'b01100011;
			9'd41:OUT=8'b01100010;
			9'd42:OUT=8'b01100010;
			9'd43:OUT=8'b01100001;
			9'd44:OUT=8'b01100000;
			9'd45:OUT=8'b01100000;
			9'd46:OUT=8'b01011111;		
			9'd47:OUT=8'b01011110;
			9'd48:OUT=8'b01011101;	
			9'd49:OUT=8'b01011101;
			9'd50:OUT=8'b01011100;
			9'd51:OUT=8'b01011011;
			9'd52:OUT=8'b01011011;
			9'd53:OUT=8'b01011010;
			9'd54:OUT=8'b01011001;
			9'd55:OUT=8'b01011000;
			9'd56:OUT=8'b01011000;
			9'd57:OUT=8'b01010111;
			9'd58:OUT=8'b01010110;
			9'd59:OUT=8'b01010110;
			9'd60:OUT=8'b01010101;
			9'd61:OUT=8'b01010100;
			9'd62:OUT=8'b01010011;
			9'd63:OUT=8'b01010011;
			9'd64:OUT=8'b01010010;
			9'd65:OUT=8'b01010001;
			9'd66:OUT=8'b01010001;
			9'd67:OUT=8'b01010000;
			9'd68:OUT=8'b01001111;
			9'd69:OUT=8'b01001110;
			9'd70:OUT=8'b01001110;
			9'd71:OUT=8'b01001101;
			9'd72:OUT=8'b01001100;
			9'd73:OUT=8'b01001100;
			9'd74:OUT=8'b01001011;
			9'd75:OUT=8'b01001010;
			9'd76:OUT=8'b01001001;
			9'd77:OUT=8'b01001001;
			9'd78:OUT=8'b01001000;
			9'd79:OUT=8'b01000111;
			9'd80:OUT=8'b01000111;
			9'd81:OUT=8'b01000110;
			9'd82:OUT=8'b01000101;
			9'd83:OUT=8'b01000100;
			9'd84:OUT=8'b01000100;
			9'd85:OUT=8'b01000011;
			9'd86:OUT=8'b01000010;
			9'd87:OUT=8'b01000010;
			9'd88:OUT=8'b01000001;
			9'd89:OUT=8'b01000000;
			9'd90:OUT=8'b01000000;
			9'd91:OUT=8'b00111111;
			9'd92:OUT=8'b00111110;
			9'd93:OUT=8'b00111101;
			9'd94:OUT=8'b00111000;
			9'd95:OUT=8'b00111100;
			9'd96:OUT=8'b00111011;
			9'd97:OUT=8'b00111011;
			9'd98:OUT=8'b00111010;
			9'd99:OUT=8'b00111001;
			9'd100:OUT=8'b00111000;
			9'd101:OUT=8'b00111000;
			9'd102:OUT=8'b00110111;
			9'd103:OUT=8'b00110110;
			9'd104:OUT=8'b00110110;
			9'd105:OUT=8'b00110101;
			9'd106:OUT=8'b00110100;
			9'd107:OUT=8'b00110011;
			9'd108:OUT=8'b00110011;
			9'd109:OUT=8'b00110010;
			9'd110:OUT=8'b00110001;
			9'd111:OUT=8'b00110001;
			9'd112:OUT=8'b00110000;
			9'd113:OUT=8'b00101111;
			9'd114:OUT=8'b00101110;
			9'd115:OUT=8'b00101110;
			9'd116:OUT=8'b00101101;
			9'd117:OUT=8'b00101100;
			9'd118:OUT=8'b00101100;
			9'd119:OUT=8'b00101011;
			9'd120:OUT=8'b00101010;
			9'd121:OUT=8'b00101001;
			9'd122:OUT=8'b00101001;
			9'd123:OUT=8'b00101000;
			9'd124:OUT=8'b00100111;
			9'd125:OUT=8'b00100111;
			9'd126:OUT=8'b00100110;
			9'd127:OUT=8'b00100101;
			9'd128:OUT=8'b00100100;
			9'd129:OUT=8'b00100100;
			9'd130:OUT=8'b00100011;
			9'd131:OUT=8'b00100010;
			9'd132:OUT=8'b00100010;
			9'd133:OUT=8'b00100001;
			9'd134:OUT=8'b00100000;
			9'd135:OUT=8'b00100000;
			9'd136:OUT=8'b00011111;
			9'd137:OUT=8'b00011110;
			9'd138:OUT=8'b00011101;
			9'd139:OUT=8'b00011101;
			9'd140:OUT=8'b00011100;
			9'd141:OUT=8'b00011011;
			9'd142:OUT=8'b00011011;
			9'd143:OUT=8'b00011010;
			9'd144:OUT=8'b00011001;
			9'd145:OUT=8'b00011000;
			9'd146:OUT=8'b00011000;
			9'd147:OUT=8'b00010111;
			9'd148:OUT=8'b00010110;
			9'd149:OUT=8'b00010110;
			9'd150:OUT=8'b00010101;
			9'd151:OUT=8'b00010100;
			9'd152:OUT=8'b00010011;
			9'd153:OUT=8'b00010011;
			9'd154:OUT=8'b00010010;
			9'd155:OUT=8'b00010001;
			9'd156:OUT=8'b00010001;
			9'd157:OUT=8'b00010000;
			9'd158:OUT=8'b00001111;
			9'd159:OUT=8'b00001110;
			9'd160:OUT=8'b00001110;
			9'd161:OUT=8'b00001101;
			9'd162:OUT=8'b00001100;
			9'd163:OUT=8'b00001100;
			9'd164:OUT=8'b00001011;
			9'd165:OUT=8'b00001010;
			9'd166:OUT=8'b00001001;
			9'd167:OUT=8'b00001001;
			9'd168:OUT=8'b00001000;
			9'd169:OUT=8'b00000111;
			9'd170:OUT=8'b00000111;
			9'd171:OUT=8'b00000110;
			9'd172:OUT=8'b00000101;
			9'd173:OUT=8'b00000100;
			9'd174:OUT=8'b00000100;
			9'd175:OUT=8'b00000011;
			9'd176:OUT=8'b00000010;
			9'd177:OUT=8'b00000010;
			9'd178:OUT=8'b00000001;
			9'd179:OUT=8'b00000000;
			9'd180:OUT=8'b00000000;
			9'd181:OUT=8'b11111111;
			9'd182:OUT=8'b11111110;
			9'd183:OUT=8'b11111101;
			9'd184:OUT=8'b11111101;
			9'd185:OUT=8'b11111100;
			9'd186:OUT=8'b11111011;
			9'd187:OUT=8'b11111011;
			9'd188:OUT=8'b11111010;
			9'd189:OUT=8'b11111001;
			9'd190:OUT=8'b11111000;
			9'd191:OUT=8'b11111000;
			9'd192:OUT=8'b11110111;
			9'd193:OUT=8'b11110110;
			9'd194:OUT=8'b11110110;
			9'd195:OUT=8'b11110101;
			9'd196:OUT=8'b11110100;
			9'd197:OUT=8'b11110011;
			9'd198:OUT=8'b11110011;
			9'd199:OUT=8'b11110010;
			9'd200:OUT=8'b11110001;
			9'd201:OUT=8'b11110001;
			9'd202:OUT=8'b11110000;
			9'd203:OUT=8'b11101111;
			9'd204:OUT=8'b11101110;
			9'd205:OUT=8'b11101110;
			9'd206:OUT=8'b11101101;
			9'd207:OUT=8'b11101100;
			9'd208:OUT=8'b11101100;
			9'd209:OUT=8'b11101011;
			9'd210:OUT=8'b11101010;
			9'd211:OUT=8'b11101001;
			9'd212:OUT=8'b11101001;
			9'd213:OUT=8'b11101000;
			9'd214:OUT=8'b11100111;
			9'd215:OUT=8'b11100111;
			9'd216:OUT=8'b11100110;
			9'd217:OUT=8'b11100101;
			9'd218:OUT=8'b11100100;
			9'd219:OUT=8'b11100100;
			9'd220:OUT=8'b11100011;
			9'd221:OUT=8'b11100010;
			9'd222:OUT=8'b11100010;
			9'd223:OUT=8'b11100001;
			9'd224:OUT=8'b11100000;
			9'd225:OUT=8'b11100000;
			9'd226:OUT=8'b11011111;
			9'd227:OUT=8'b11011110;
			9'd228:OUT=8'b11011101;
			9'd229:OUT=8'b11011101;
			9'd230:OUT=8'b11011100;
			9'd231:OUT=8'b11011011;
			9'd232:OUT=8'b11011011;
			9'd233:OUT=8'b11011010;
			9'd234:OUT=8'b11011001;
			9'd235:OUT=8'b11011000;
			9'd236:OUT=8'b11011000;
			9'd237:OUT=8'b11010111;
			9'd238:OUT=8'b11010110;
			9'd239:OUT=8'b11010110;
			9'd240:OUT=8'b11010101;
			9'd241:OUT=8'b11010100;
			9'd242:OUT=8'b11010011;
			9'd243:OUT=8'b11010011;
			9'd244:OUT=8'b11010010;
			9'd245:OUT=8'b11010001;
			9'd246:OUT=8'b11010001;
			9'd247:OUT=8'b11010000;
			9'd248:OUT=8'b11001111;
			9'd249:OUT=8'b11001110;
			9'd250:OUT=8'b11001110;
			9'd251:OUT=8'b11001101;
			9'd252:OUT=8'b11001100;
			9'd253:OUT=8'b11001100;
			9'd254:OUT=8'b11001011;
			9'd255:OUT=8'b11001010;
			9'd256:OUT=8'b11001001;
			9'd257:OUT=8'b11001001;
			9'd258:OUT=8'b11001000;
			9'd259:OUT=8'b11000111;
			9'd260:OUT=8'b11000111;
			9'd261:OUT=8'b11000110;
			9'd262:OUT=8'b11000101;
			9'd263:OUT=8'b11000100;
			9'd264:OUT=8'b11000100;
			9'd265:OUT=8'b11000011;
			9'd266:OUT=8'b11000010;
			9'd267:OUT=8'b11000010;
			9'd268:OUT=8'b11000001;
			9'd269:OUT=8'b11000000;
			9'd270:OUT=8'b11000000;
			9'd271:OUT=8'b10111111;
			9'd272:OUT=8'b10111110;
			9'd273:OUT=8'b10111101;
			9'd274:OUT=8'b10111101;
			9'd275:OUT=8'b10111100;
			9'd276:OUT=8'b10111011;
			9'd277:OUT=8'b10111011;
			9'd278:OUT=8'b10111010;
			9'd279:OUT=8'b10111001;
			9'd280:OUT=8'b10111000;
			9'd281:OUT=8'b10111000;
			9'd282:OUT=8'b10110111;
			9'd283:OUT=8'b10110110;
			9'd284:OUT=8'b10110110;
			9'd285:OUT=8'b10110101;
			9'd286:OUT=8'b10110100;
			9'd287:OUT=8'b10110011;
			9'd288:OUT=8'b10110011;
			9'd289:OUT=8'b10110010;
			9'd290:OUT=8'b10110001;
			9'd291:OUT=8'b10110001;
			9'd292:OUT=8'b10110000;
			9'd293:OUT=8'b10101111;
			9'd294:OUT=8'b10101110;
			9'd295:OUT=8'b10101110;
			9'd296:OUT=8'b10101101;
			9'd297:OUT=8'b10101100;
			9'd298:OUT=8'b10101100;
			9'd299:OUT=8'b10101011;
			9'd300:OUT=8'b10101010;
			9'd301:OUT=8'b10101001;
			9'd302:OUT=8'b10101001;
			9'd303:OUT=8'b10101000;
			9'd304:OUT=8'b10100111;
			9'd305:OUT=8'b10100111;
			9'd306:OUT=8'b10100110;
			9'd307:OUT=8'b10100101;
			9'd308:OUT=8'b10100100;
			9'd309:OUT=8'b10100100;
			9'd310:OUT=8'b10100011;
			9'd311:OUT=8'b10100010;
			9'd312:OUT=8'b10100010;
			9'd313:OUT=8'b10100001;
			9'd314:OUT=8'b10100000;
			9'd315:OUT=8'b10100000;
			9'd316:OUT=8'b10011111;
			9'd317:OUT=8'b10011110;
			9'd318:OUT=8'b10011101;
			9'd319:OUT=8'b10011101;
			9'd320:OUT=8'b10011100;
			9'd321:OUT=8'b10011011;
			9'd322:OUT=8'b10011011;
			9'd323:OUT=8'b10011010;
			9'd324:OUT=8'b10011001;
			9'd325:OUT=8'b10011000;
			9'd326:OUT=8'b10011000;
			9'd327:OUT=8'b10010111;
			9'd328:OUT=8'b10010110;
			9'd329:OUT=8'b10010110;
			9'd330:OUT=8'b10010101;
			9'd331:OUT=8'b10010100;
			9'd332:OUT=8'b10010011;
			9'd333:OUT=8'b10010011;
			9'd334:OUT=8'b10010010;
			9'd335:OUT=8'b10010001;
			9'd336:OUT=8'b10010001;
			9'd337:OUT=8'b10010000;
			9'd338:OUT=8'b10001111;
			9'd339:OUT=8'b10001110;
			9'd340:OUT=8'b10001110;

			default OUT=8'b00000000;
		endcase



endmodule
